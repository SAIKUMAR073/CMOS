***Write Operation
VDD 3 0 dc 5V
Vbit 5 0 dc 5V
Vbitb 6 0 dc 0V
Vw 4 0 pulse(5 0 0 0 0 50ms 100ms)
C1 5 0 0.1p
C2 6 0 0.1
.model nmod nmos level = 54 version = 4.7
.model pmod pmos level = 54 version = 4.7
M1 1 2 3 3 pmod w = 100u l = 10u
M2 1 2 0 0 nmod w = 100u l = 10u
M3 2 1 3 3 pmod w = 100u l = 10u
M4 2 1 0 0 nmod w = 100u l = 10u
M5 1 4 5 0 nmod w = 100u l = 10u
M6 2 4 6 0 nmod w = 100u l = 10u
.tran 0.01ms 200ms 
.control
run
plot V(4)
plot V(1)
plot V(2)
.endc
.end